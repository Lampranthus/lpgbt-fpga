library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity prbs7_64b_generator is
    generic(
        INIT_c                  : in std_logic_vector(63 downto 0)
    );
    port (
        reset_i          : in  std_logic;
        clk_i            : in  std_logic;
        clk_enable_i     : in  std_logic;

        prbs_word_o      : out std_logic_vector(63 downto 0);
        rdy_o            : out std_logic
    );
end prbs7_64b_generator;

architecture rtl of prbs7_64b_generator is
    signal feedback_reg         : std_logic_vector(63 downto 0) := INIT_c;
    signal prbs_word_s          : std_logic_vector(63 downto 0) := INIT_c;

begin

    -- PRBS7 equation: x^7 + x^6 + 1
    -- LSB first

    prbs7_proc: process(reset_i, clk_i)
    begin

        if reset_i = '1' then
            feedback_reg <= INIT_c;
            prbs_word_s  <= INIT_c;
            rdy_o        <= '0';

        elsif rising_edge(clk_i) then

            if clk_enable_i = '1' then

                prbs_word_s  <= feedback_reg;
                rdy_o        <= '1';

                feedback_reg(0) <= feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2);
                feedback_reg(1) <= feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3);
                feedback_reg(2) <= feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4);
                feedback_reg(3) <= feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5);
                feedback_reg(4) <= feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0);
                feedback_reg(5) <= feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1);
                feedback_reg(6) <= feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2);
                feedback_reg(7) <= feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3);
                feedback_reg(8) <= feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4);
                feedback_reg(9) <= feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5);
                feedback_reg(10) <= feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0);
                feedback_reg(11) <= feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1);
                feedback_reg(12) <= feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2);
                feedback_reg(13) <= feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3);
                feedback_reg(14) <= feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4);
                feedback_reg(15) <= feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5);
                feedback_reg(16) <= feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0);
                feedback_reg(17) <= feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1);
                feedback_reg(18) <= feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2);
                feedback_reg(19) <= feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3);
                feedback_reg(20) <= feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4);
                feedback_reg(21) <= feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5);
                feedback_reg(22) <= feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0);
                feedback_reg(23) <= feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1);
                feedback_reg(24) <= feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2);
                feedback_reg(25) <= feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3);
                feedback_reg(26) <= feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4);
                feedback_reg(27) <= feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5);
                feedback_reg(28) <= feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0);
                feedback_reg(29) <= feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1);
                feedback_reg(30) <= feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2);
                feedback_reg(31) <= feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3);
                feedback_reg(32) <= feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4);
                feedback_reg(33) <= feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5);
                feedback_reg(34) <= feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0);
                feedback_reg(35) <= feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1);
                feedback_reg(36) <= feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2);
                feedback_reg(37) <= feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3);
                feedback_reg(38) <= feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4);
                feedback_reg(39) <= feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5);
                feedback_reg(40) <= feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0);
                feedback_reg(41) <= feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1);
                feedback_reg(42) <= feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2);
                feedback_reg(43) <= feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3);
                feedback_reg(44) <= feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4);
                feedback_reg(45) <= feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5);
                feedback_reg(46) <= feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0);
                feedback_reg(47) <= feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1);
                feedback_reg(48) <= feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2);
                feedback_reg(49) <= feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3);
                feedback_reg(50) <= feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4);
                feedback_reg(51) <= feedback_reg(1) xor feedback_reg(0) xor feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5);
                feedback_reg(52) <= feedback_reg(2) xor feedback_reg(1) xor feedback_reg(1) xor feedback_reg(0);
                feedback_reg(53) <= feedback_reg(3) xor feedback_reg(2) xor feedback_reg(2) xor feedback_reg(1);
                feedback_reg(54) <= feedback_reg(4) xor feedback_reg(3) xor feedback_reg(3) xor feedback_reg(2);
                feedback_reg(55) <= feedback_reg(5) xor feedback_reg(4) xor feedback_reg(4) xor feedback_reg(3);
                feedback_reg(56) <= feedback_reg(6) xor feedback_reg(5) xor feedback_reg(5) xor feedback_reg(4);
                feedback_reg(57) <= feedback_reg(0) xor feedback_reg(6) xor feedback_reg(5);
                feedback_reg(58) <= feedback_reg(1) xor feedback_reg(0);
                feedback_reg(59) <= feedback_reg(2) xor feedback_reg(1);
                feedback_reg(60) <= feedback_reg(3) xor feedback_reg(2);
                feedback_reg(61) <= feedback_reg(4) xor feedback_reg(3);
                feedback_reg(62) <= feedback_reg(5) xor feedback_reg(4);
                feedback_reg(63) <= feedback_reg(6) xor feedback_reg(5);

            end if;

        end if;

    end process;

    prbs_word_o   <= prbs_word_s;

end rtl;
